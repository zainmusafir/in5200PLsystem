
package kb_axi4stream_typedef_pkg;

   typedef enum {TX, RX, TXRX, NOP} axi4stream_transaction_type_t;
    
endpackage: kb_axi4stream_typedef_pkg

