package psif_odi_spi_pkg;
   
   import uvm_pkg::*;

   import tb_env_pkg::*;
   import base_test_pkg::*;
   import base_seq_pkg::*;
   import axi4params_pkg::*;
 
   `include "uvm_macros.svh";
   `include "psif_odi_spi_seq.svh";
   `include "psif_odi_spi_seq_virtual.svh";
   `include "psif_odi_spi_test.svh";
  
endpackage // psif_odi_spi_pkg
   
