package psif_aui_aurora_pkg;
   
   import uvm_pkg::*;

//   import interrupt_handler_pkg::*;
   import tb_env_pkg::*;
   import tb_env_base_pkg::*;
   import base_test_pkg::*;
   import base_seq_pkg::*;
   import kb_axi4stream_agent_pkg::*; 

   import probe_pkg::*;
  
   `include "uvm_macros.svh";

   import axi4params_pkg::*;  

   `include "aurora_seq.svh";
   `include "psif_aui_aurora_init_seq.svh";
   `include "psif_aui_aurora_loop_seq.svh";
   `include "psif_aui_aurora_tx_seq.svh";
   `include "psif_aui_aurora_rx_seq.svh";
   `include "psif_aui_aurora_seq_virtual.svh";
   `include "psif_aui_aurora_test.svh";
  
endpackage // psif_aui_aurora_pkg
   
