package psif_ram_pkg;
   
   import uvm_pkg::*;

   import tb_env_pkg::*;
   import base_test_pkg::*;
   import base_seq_pkg::*;
   import axi4params_pkg::*;
   
   `include "uvm_macros.svh";
   `include "psif_ram_test.svh";
  
endpackage // psif_ram_pkg
   
