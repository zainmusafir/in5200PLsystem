

interface reset_agent_if(input clk);

   logic  rst;
      
endinterface // reset_agent_if

