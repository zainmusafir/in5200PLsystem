--
-- Written by Ryan Kim, Digilent Inc.
-- Modified by Michael Mattioli
--
-- Description: Top level controller that controls the OLED display.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity oled_ctrl is
    generic (
      SIMULATION_MODE : string);
    port (  clk           : in  std_logic;
            rst           : in  std_logic;
            oledbyte3_0   : in  std_logic_vector(31 downto 0);
            oledbyte7_4   : in  std_logic_vector(31 downto 0);
            oledbyte11_8  : in  std_logic_vector(31 downto 0);
            oledbyte15_12 : in  std_logic_vector(31 downto 0);  
            oled_sdin     : out std_logic;
            oled_sclk     : out std_logic;
            oled_dc       : out std_logic;
            oled_res      : out std_logic;
            oled_vbat     : out std_logic;
            oled_vdd      : out std_logic);
end oled_ctrl;

architecture behavioral of oled_ctrl is

    component oled_init is
        generic (
          SIMULATION_MODE : string);
        port (  clk         : in std_logic;
                rst         : in std_logic;
                en          : in std_logic;
                sdout       : out std_logic;
                oled_sclk   : out std_logic;
                oled_dc     : out std_logic;
                oled_res    : out std_logic;
                oled_vbat   : out std_logic;
                oled_vdd    : out std_logic;
                fin         : out std_logic);
    end component;

    component oled_ex is
        generic (
          SIMULATION_MODE : string);
        port (  clk           : in  std_logic;
                rst           : in  std_logic;
                en            : in  std_logic;
                line1_1       : in  string;
                line3_1       : in  string;
                line1_2       : in  string;
                oledbyte3_0   : in  std_logic_vector(31 downto 0);
                oledbyte7_4   : in  std_logic_vector(31 downto 0);
                oledbyte11_8  : in  std_logic_vector(31 downto 0);
                oledbyte15_12 : in  std_logic_vector(31 downto 0);
                sdout         : out std_logic;
                oled_sclk     : out std_logic;
                oled_dc       : out std_logic;
                fin           : out std_logic;
                alphabet_done_str : out std_logic); -- ADDED alphabet_done strobe signal for simulation/testbench purposes

    end component;

    type states is (Idle, OledInitialize, OledExample, Done);

    signal current_state : states := Idle;

    signal init_en          : std_logic := '0';
    signal init_done        : std_logic;
    signal init_sdata       : std_logic;
    signal init_spi_clk     : std_logic;
    signal init_dc          : std_logic;

    signal example_en       : std_logic := '0';
    signal example_sdata    : std_logic;
    signal example_spi_clk  : std_logic;
    signal example_dc       : std_logic;
    signal example_done     : std_logic;

    signal alphabet_done_str : std_logic; -- ADDED alphabet_done strobe signal for simulation/testbench purposes

    constant line1_1 : string(1 to 16):= "Welcome:        ";
    constant line3_1 : string(1 to 16):= "  IN5200 lab    ";    
    constant line1_2 : string(1 to 16):= "Lab output:     ";
    
begin

    Initialize: oled_init
      generic map (
        SIMULATION_MODE => SIMULATION_MODE)
      port map (clk,
                rst,
                init_en,
                init_sdata,
                init_spi_clk,
                init_dc,
                oled_res,
                oled_vbat,
                oled_vdd,
                init_done);

    Example: oled_ex
      generic map (
        SIMULATION_MODE => SIMULATION_MODE)
      port map ( clk,
                 rst,
                 example_en,
                 line1_1,
                 line3_1,
                 line1_2,
                 oledbyte3_0,   
                 oledbyte7_4,   
                 oledbyte11_8,  
                 oledbyte15_12,
                 example_sdata,
                 example_spi_clk,
                 example_dc,
                 example_done,
                 alphabet_done_str); -- ADDED alphabet_done strobe signal for simulation/testbench purposes

    -- MUXes to indicate which outputs are routed out depending on which block is enabled
    oled_sdin <= init_sdata when current_state = OledInitialize else example_sdata;
    oled_sclk <= init_spi_clk when current_state = OledInitialize else example_spi_clk;
    oled_dc <= init_dc when current_state = OledInitialize else example_dc;
    -- End output MUXes

    -- MUXes that enable blocks when in the proper states
    init_en <= '1' when current_state = OledInitialize else '0';
    example_en <= '1' when current_state = OledExample else '0';
    -- End enable MUXes

    process (clk)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                current_state <= Idle;
            else
                case current_state is
                    when Idle =>
                        current_state <= OledInitialize;
                    -- Go through the initialization sequence
                    when OledInitialize =>
                        if init_done = '1' then
                            current_state <= OledExample;
                        end if;
                    -- Do example and do nothing when finished
                    when OledExample =>
                        if example_done = '1' then
                            current_state <= Done;
                        end if;
                    -- Do nthing
                    when Done =>
                        current_state <= Done;
                    when others =>
                        current_state <= Idle;
                end case;
            end if;
        end if;
    end process;

end behavioral;
