package psif_scu_pkg;
   
   import uvm_pkg::*;

   import tb_env_pkg::*;
   import base_test_pkg::*;
   import base_seq_pkg::*;
   import axi4params_pkg::*;
 
   `include "uvm_macros.svh";
   `include "psif_scu_seq.svh";
   `include "psif_scu_seq_virtual.svh";
   `include "psif_scu_test.svh";
  
endpackage // psif_scu_pkg
   