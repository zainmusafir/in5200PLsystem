
//----------------------------------------------------------------------
// oled_spi_agent
//----------------------------------------------------------------------
class oled_spi_agent extends uvm_agent;

  // factory registration macro
  `uvm_component_utils(oled_spi_agent)   

  // configuration object
  oled_spi_agent_config m_cfg;

  // internal components
  oled_spi_agent_driver   m_driver;
  oled_spi_agent_monitor  m_monitor;
  uvm_sequencer #(oled_spi_agent_item) sequencer;

  //--------------------------------------------------------------------
  // new
  //--------------------------------------------------------------------
  function new(string name = "oled_spi_agent", 
               uvm_component parent = null);
    super.new(name, parent);
  endfunction: new

  //--------------------------------------------------------------------
  // build_phase
  //--------------------------------------------------------------------
  virtual function void build_phase(uvm_phase phase);
    
    if(!uvm_config_db #(oled_spi_agent_config)::get(this, "", "oled_spi_agent_config", m_cfg)) begin
      `uvm_error("build_phase", "oled_spi_agent_config not found")
    end    

    m_monitor   = oled_spi_agent_monitor::type_id::create("m_monitor",this);
   
    // Driver and Sequencer only built if agent is active
    if (m_cfg.is_active == UVM_ACTIVE) begin
      m_driver   = oled_spi_agent_driver::type_id::create("m_driver",this);
      sequencer  = uvm_sequencer #(oled_spi_agent_item)::type_id::create("sequencer",this); 
      m_cfg.sequencer=sequencer;
    end 
  endfunction: build_phase

  //--------------------------------------------------------------------
  // connect_phase
  //--------------------------------------------------------------------
  virtual function void connect_phase(uvm_phase phase);

    // Monitor is always connected
//    m_monitor.ap.connect(ap);
    m_monitor.m_cfg = m_cfg;
    
    // Driver and Sequencer only connected if agent is active    
    if (m_cfg.is_active == UVM_ACTIVE) begin
      m_driver.m_cfg=m_cfg; // The virtual interface is included in the m_cfg class!!!
      m_driver.seq_item_port.connect(sequencer.seq_item_export);   
    end     
    
  endfunction: connect_phase

endclass: oled_spi_agent

