

interface oled_spi_agent_if(input clk);

   logic oled_sdin;
   logic oled_sclk;
   logic oled_dc;
   logic oled_res;
   logic oled_vbat;
   logic oled_vdd;
      
endinterface // oled_spi_agent_if

