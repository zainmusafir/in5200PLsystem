   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(1))   aes_inv_cipher_probe_ap_clk(ap_clk);
   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(1))   aes_inv_cipher_probe_bypass(bypass);
   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(1))   aes_inv_cipher_probe_ap_start(ap_start);
   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(1))   aes_inv_cipher_probe_ap_done(ap_done);
   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(8))   aes_inv_cipher_probe_out_r_tdata(out_r_tdata);
   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(1))   aes_inv_cipher_probe_out_r_tvalid(out_r_tvalid);
   bind aes_inv_cipher : tb_top.mla_top.mla_pl.zu_0.aes128_inv_cipher_0   probe_itf #(.WIDTH(1))   aes_inv_cipher_probe_out_r_tready(out_r_tready);
